class driver;

  virtual uart_if vif;
  transaction tr;

  mailbox #(transaction) mbx;
  mailbox #(bit [7:0]) mbxds;

  event drvnext;

  bit [7:0] din;
  bit wr = 0;
  bit [7:0] datarx;

  function new(mailbox #(bit [7:0]) mbxds,
               mailbox #(transaction) mbx);
    this.mbx   = mbx;
    this.mbxds = mbxds;
  endfunction

  task reset();
    vif.rst   <= 1'b1;
    vif.dintx <= 0;
    vif.newd  <= 0;
    vif.rx    <= 1'b1;

    repeat(5) @(posedge vif.uclktx);
    vif.rst <= 1'b0;
    @(posedge vif.uclktx);

    $display("[DRV] : RESET DONE");
    $display("----------------------------------------");
  endtask

  task run();
    forever begin
      mbx.get(tr);

      // WRITE OPERATION
      if(tr.oper == 1'b0) begin
        @(posedge vif.uclktx);
        vif.rst  <= 1'b0;
        vif.newd <= 1'b1;
        vif.rx   <= 1'b1;
        vif.dintx = tr.dintx;

        @(posedge vif.uclktx);
        vif.newd <= 1'b0;

        mbxds.put(tr.dintx);
        $display("[DRV]: Data Sent : %0d", tr.dintx);

        wait(vif.donetx == 1'b1);
        ->drvnext;
      end

      // READ OPERATION
      else begin
        @(posedge vif.uclkrx);
        vif.rst  <= 1'b0;
        vif.rx   <= 1'b0;
        vif.newd <= 1'b0;

        @(posedge vif.uclkrx);

        for(int i = 0; i <= 7; i++) begin
          @(posedge vif.uclkrx);
          vif.rx = $urandom;
          datarx[i] = vif.rx;
        end

        mbxds.put(datarx);
        $display("[DRV]: Data RCVD : %0d", datarx);

        wait(vif.donerx == 1'b1);
        vif.rx <= 1'b1;

        ->drvnext;
      end
    end
  endtask

endclass
